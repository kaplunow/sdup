module cordic_beh_fixedpoint();
//12:10 data representation
parameter real FXP_SCALE = 1024.0; //scale factor = 2^10
parameter integer FXP_SCALE_SHIFT = 10;
/**
* Cordic algorithm
*/
reg signed [11:0] t_angle = 0.8 * FXP_SCALE; //Input angle

//Table of arctan (1/2^i)
// Note. Table initialization below is not correct for Verilog. Select System-Verilog mode
// in your simulator in the case of syntax errors
reg signed [11:0] arctan[0:10];
reg signed [11:0] Kn = 0.607252937 * FXP_SCALE; //Cordic scaling factor for 10 iterationsreg signed [11:0] Kn = 0.607252937 * FXP_SCALE;
//Variables
reg signed [11:0] cos = 1.0 * FXP_SCALE; //Initial condition
reg signed [11:0] sin = 0.0 * FXP_SCALE;

reg signed [11:0] angle = 0.0 * FXP_SCALE; //Running angle

reg signed [23:0] Kn_sin;
reg signed [23:0] Kn_cos;
integer i;
reg signed [11:0] tmp;

initial //Execute only once
begin
    //FXP_SCALED atan values, generated by python script
	arctan[0]  = 804;
	arctan[1]  = 475;
	arctan[2]  = 251;
	arctan[3]  = 127;
	arctan[4]  = 64;
	arctan[5]  = 32;
	arctan[6]  = 16;
	arctan[7]  = 8;
	arctan[8]  = 4;
	arctan[9]  = 2;
	arctan[10] = 1;

	for ( i = 0; i < 11; i = i + 1) //Ten algorithm iterations
	begin
		if( t_angle > angle )
		begin
			angle = angle + arctan[i];
			tmp = cos - ( sin >>> i );
			sin = ( cos >>> i ) + sin;
			cos = tmp;
		end
		else
		begin
			angle = angle - arctan[i];
			tmp = cos + ( sin >>> i );
			sin = - ( cos >>> i) + sin;
			cos = tmp;
		end //if
	end //for
	//Scale sin/cos values
	Kn_sin = Kn * sin;
	sin = Kn_sin >>> FXP_SCALE_SHIFT;
	Kn_cos = Kn * cos;
	cos = Kn_cos >>> FXP_SCALE_SHIFT;
	
	$display("sin=%f, cos=%f", sin/FXP_SCALE, cos/FXP_SCALE);
end
    
endmodule
